package shared_pkg;

    bit test_finished;
    int error_count, correct_count;   
endpackage
